library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity datapath is
    port (
        clk, clr, ld_floor, ld_call : in  bit;
        
        -- chaves dos MUXs, que vem do controlador:
        ctrl_s1, ctrl_s0 : in bit;

        -- andar que o elevador foi chamado 
        call_floor_in : in  BIT_VECTOR(1 downto 0);

        -- flags para o controlador 
        lt, eq, gt : out bit;

        -- saida para display / monitoramento
        display_floor : out BIT_VECTOR(1 downto 0)
    );
end entity datapath;

architecture rtl of datapath is
    component reg2 is
        port (
            clk : in bit;
            ld  : in bit;
            clr : in bit;
            d   : in BIT_VECTOR(1 downto 0);
            q   : out BIT_VECTOR(1 downto 0)
        );
    end component;

    component Mux4x1 is
        port (
            i3, i2, i1, i0 : in bit;
            s1, s0         : in bit;
            d              : out bit
        );
    end component;

    component comparador_2bits is
        port (
            b1, b0, a1, a0: in bit;
            l_t, e_t, g_t : out bit
        );
    end component;

    component subtrator_2bits is
        port (
            a0, a1, b0, b1 : in bit;
            s0, s1, co     : out bit
        );
    end component;

    component somador_2bits is
        port (
            a0, a1, b0, b1 : in bit;
            s0, s1, co     : out bit
        );
    end component;

    -- sinais internos (2 bits)
    signal r_current     : BIT_VECTOR(1 downto 0);
    signal r_call_floor  : BIT_VECTOR(1 downto 0);
    signal r_next        : BIT_VECTOR(1 downto 0);
    signal r_sum         : BIT_VECTOR(1 downto 0);
    signal r_sub         : BIT_VECTOR(1 downto 0);

    -- saidas pro comparador
    signal comp_lt, comp_eq, comp_gt : bit;

    -- carry outs (nao usados)
    signal co_sum, co_sub : bit;

begin
    -- registrador do andar atual
    reg_current : reg2
        port map(
            clk => clk,
            ld  => ld_floor,
            clr => clr,
            d   => r_next,
            q   => r_current
        );

    -- registrador do andar chamado
    reg_call_floor : reg2
        port map(
            clk => clk,
            ld  => ld_call,    
            clr => clr,
            d   => call_floor_in,
            q   => r_call_floor
        );

    -- comparacao entre current_floor e call_floor
    comp : comparador_2bits
        port map(
            b1 => r_current(1),
            b0 => r_current(0),
            a1 => r_call_floor(1),
            a0 => r_call_floor(0),
            l_t => comp_lt,
            e_t => comp_eq,
            g_t => comp_gt
        );

    lt <= comp_lt;
    eq <= comp_eq;
    gt <= comp_gt;

    -- soma com 1
    somador_unitario : somador_2bits
        port map(
            a0 => r_current(0),
            a1 => r_current(1),
            b0 => '1',
            b1 => '0',
            s0 => r_sum(0),
            s1 => r_sum(1),
            co => co_sum
        );

    -- subtrai com 1
    subtrator_unitario : subtrator_2bits
        port map(
            a0 => r_current(0),
            a1 => r_current(1),
            b0 => '1',
            b1 => '0',
            s0 => r_sub(0),
            s1 => r_sub(1),
            co => co_sub
        );

    ------------------------------------------------------------------------
    -- Mux 4x1 (implementado por 2 instancias, 1 bit por vez)
    -- selecao: s1 = comp_gt, s0 = comp_lt
    -- codificacao usada:
    --   s1 s0 = 00 -> i0 = manter (r_current)
    --   s1 s0 = 01 -> i1 = descer (r_sub)
    --   s1 s0 = 10 -> i2 = subir  (r_sum)
    --   s1 s0 = 11 -> i3 = manter (r_current)
    ------------------------------------------------------------------------
    mux_output_0 : Mux4x1
        port map(
            i3 => r_current(0),
            i2 => r_sum(0),
            i1 => r_sub(0),
            i0 => r_current(0),
            s1 => ctrl_s1,
            s0 => ctrl_s0,
            d  => r_next(0)
        );

    mux_output_1 : Mux4x1
        port map(
            i3 => r_current(1),
            i2 => r_sum(1),
            i1 => r_sub(1),
            i0 => r_current(1),
            s1 => ctrl_s1,
            s0 => ctrl_s0,
            d  => r_next(1)
        );

    display_floor <= r_current;

end architecture rtl;
